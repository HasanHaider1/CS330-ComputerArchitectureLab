module tb2
(

);